hello verifworks
